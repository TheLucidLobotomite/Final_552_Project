module decode (
    
) (
    ports
);
    
endmodule
module ExtoMEM();

endmodule
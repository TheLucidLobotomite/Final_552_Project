module hart #(
    // After reset, the program counter (PC) should be initialized to this
    // address and start executing instructions from there.
    parameter RESET_ADDR = 32'h00000000
) (
    // Global clock.
    input  wire        i_clk,
    // Synchronous active-high reset.
    input  wire        i_rst,
    // Instruction fetch goes through a read only instruction memory (imem)
    // port. The port accepts a 32-bit address (e.g. from the program counter)
    // per cycle and combinationally returns a 32-bit instruction word. This
    // is not representative of a realistic memory interface; it has been
    // modeled as more similar to a DFF or SRAM to simplify phase 3. In
    // later phases, you will replace this with a more realistic memory.
    //
    // 32-bit read address for the instruction memory. This is expected to be
    // 4 byte aligned - that is, the two LSBs should be zero.
    output wire [31:0] o_imem_raddr,
    // Instruction word fetched from memory, available on the same cycle.
    input  wire [31:0] i_imem_rdata,
    // Data memory accesses go through a separate read/write data memory (dmem)
    // that is shared between read (load) and write (stored). The port accepts
    // a 32-bit address, read or write enable, and mask (explained below) each
    // cycle. Reads are combinational - values are available immediately after
    // updating the address and asserting read enable. Writes occur on (and
    // are visible at) the next clock edge.
    //
    // Read/write address for the data memory. This should be 32-bit aligned
    // (i.e. the two LSB should be zero). See `o_dmem_mask` for how to perform
    // half-word and byte accesses at unaligned addresses.
    output wire [31:0] o_dmem_addr,
    // When asserted, the memory will perform a read at the aligned address
    // specified by `i_addr` and return the 32-bit word at that address
    // immediately (i.e. combinationally). It is illegal to assert this and
    // `o_dmem_wen` on the same cycle.
    output wire        o_dmem_ren,
    // When asserted, the memory will perform a write to the aligned address
    // `o_dmem_addr`. When asserted, the memory will write the bytes in
    // `o_dmem_wdata` (specified by the mask) to memory at the specified
    // address on the next rising clock edge. It is illegal to assert this and
    // `o_dmem_ren` on the same cycle.
    output wire        o_dmem_wen,
    // The 32-bit word to write to memory when `o_dmem_wen` is asserted. When
    // write enable is asserted, the byte lanes specified by the mask will be
    // written to the memory word at the aligned address at the next rising
    // clock edge. The other byte lanes of the word will be unaffected.
    output wire [31:0] o_dmem_wdata,
    // The dmem interface expects word (32 bit) aligned addresses. However,
    // WISC-25 supports byte and half-word loads and stores at unaligned and
    // 16-bit aligned addresses, respectively. To support this, the access
    // mask specifies which bytes within the 32-bit word are actually read
    // from or written to memory.
    //
    // To perform a half-word read at address 0x00001002, align `o_dmem_addr`
    // to 0x00001000, assert `o_dmem_ren`, and set the mask to 0b1100 to
    // indicate that only the upper two bytes should be read. Only the upper
    // two bytes of `i_dmem_rdata` can be assumed to have valid data; to
    // calculate the final value of the `lh[u]` instruction, shift the rdata
    // word right by 16 bits and sign/zero extend as appropriate.
    //
    // To perform a byte write at address 0x00002003, align `o_dmem_addr` to
    // `0x00002000`, assert `o_dmem_wen`, and set the mask to 0b1000 to
    // indicate that only the upper byte should be written. On the next clock
    // cycle, the upper byte of `o_dmem_wdata` will be written to memory, with
    // the other three bytes of the aligned word unaffected. Remember to shift
    // the value of the `sb` instruction left by 24 bits to place it in the
    // appropriate byte lane.
    output wire [ 3:0] o_dmem_mask,
    // The 32-bit word read from data memory. When `o_dmem_ren` is asserted,
    // this will immediately reflect the contents of memory at the specified
    // address, for the bytes enabled by the mask. When read enable is not
    // asserted, or for bytes not set in the mask, the value is undefined.
    input  wire [31:0] i_dmem_rdata,
	// The output `retire` interface is used to signal to the testbench that
    // the CPU has completed and retired an instruction. A single cycle
    // implementation will assert this every cycle; however, a pipelined
    // implementation that needs to stall (due to internal hazards or waiting
    // on memory accesses) will not assert the signal on cycles where the
    // instruction in the writeback stage is not retiring.
    //
    // Asserted when an instruction is being retired this cycle. If this is
    // not asserted, the other retire signals are ignored and may be left invalid.
    output wire        o_retire_valid,
    // The 32 bit instruction word of the instrution being retired. This
    // should be the unmodified instruction word fetched from instruction
    // memory.
    output wire [31:0] o_retire_inst,
    // Asserted if the instruction produced a trap, due to an illegal
    // instruction, unaligned data memory access, or unaligned instruction
    // address on a taken branch or jump.
    output wire        o_retire_trap,
    // Asserted if the instruction is an `ebreak` instruction used to halt the
    // processor. This is used for debugging and testing purposes to end
    // a program.
    output wire        o_retire_halt,
    // The first register address read by the instruction being retired. If
    // the instruction does not read from a register (like `lui`), this
    // should be 5'd0.
    output wire [ 4:0] o_retire_rs1_raddr,
    // The second register address read by the instruction being retired. If
    // the instruction does not read from a second register (like `addi`), this
    // should be 5'd0.
    output wire [ 4:0] o_retire_rs2_raddr,
    // The first source register data read from the register file (in the
    // decode stage) for the instruction being retired. If rs1 is 5'd0, this
    // should also be 32'd0.
    output wire [31:0] o_retire_rs1_rdata,
    // The second source register data read from the register file (in the
    // decode stage) for the instruction being retired. If rs2 is 5'd0, this
    // should also be 32'd0.
    output wire [31:0] o_retire_rs2_rdata,
    // The destination register address written by the instruction being
    // retired. If the instruction does not write to a register (like `sw`),
    // this should be 5'd0.
    output wire [ 4:0] o_retire_rd_waddr,
    // The destination register data written to the register file in the
    // writeback stage by this instruction. If rd is 5'd0, this field is
    // ignored and can be treated as a don't care.
    output wire [31:0] o_retire_rd_wdata,
    // The current program counter of the instruction being retired - i.e.
    // the instruction memory address that the instruction was fetched from.
    output wire [31:0] o_retire_pc,
    // the next program counter after the instruction is retired. For most
    // instructions, this is `o_retire_pc + 4`, but must be the branch or jump
    // target for *taken* branches and jumps.
    output wire [31:0] o_retire_next_pc

`ifdef RISCV_FORMAL
    ,`RVFI_OUTPUTS,
`endif
);
    /////////////////////////////////////
    // PC/Instruction Fetch Phase
    /////////////////////////////////////
    reg  [31:0] pc_reg;
    wire [31:0] pc_next;
    wire [31:0] instruction;
    wire [31:0] pc_plus_4 = pc_reg + 32'd4; //added in order to pipeline throughout
    
    assign o_imem_raddr = pc_reg;
    assign instruction = i_imem_rdata;

    always @(posedge i_clk) begin
        if (i_rst)
            pc_reg <= RESET_ADDR;
        else
            pc_reg <= pc_next;
    end
   

    /////////////////////////////////////
    // Decode Phase
    /////////////////////////////////////
    wire [31:0] o_rs1_rdata, o_rs2_rdata, o_immediate;
    wire        jump, jalr, branch;
    wire [2:0]  branch_type, i_opsel;
    wire [1:0]  rd_dest_select;
    wire [2:0]  store_sel, load_sel;
    wire        dmem_ren, dmem_wen;
    wire        i_sub, i_unsigned, i_arith, auipc, i_alu_src, i_rd_wen;
    wire [5:0]  i_format;
    wire [31:0] writeback_mux_out;

    decode iDUT_decode (
        .clk                (i_clk),
        .rst                (i_rst),
        .i_imem_rdata       (instruction),
        .writeback_mux_out  (writeback_mux_out),
        .o_rs1_data_in      (o_rs1_rdata),
        .o_rs2_data_in      (o_rs2_rdata),
        .o_immediate        (o_immediate),
        .jump               (jump),
        .jalr               (jalr),
        .branch             (branch),
        .branch_type        (branch_type),
        .rd_dest_select     (rd_dest_select),
        .store_sel          (store_sel),
        .load_sel           (load_sel),
        .o_dmem_ren         (dmem_ren),
        .o_dmem_wen         (dmem_wen),
        .i_opsel            (i_opsel),
        .i_arith            (i_arith),
        .i_unsigned         (i_unsigned),
        .i_sub              (i_sub),
        .auipc              (auipc),
        .i_alu_src          (i_alu_src),
        .i_rd_wen           (i_rd_wen),
        .i_format           (i_format)
    );

    /////////////////////////////////////
    // Execute Phase
    /////////////////////////////////////
    wire [31:0] alu_result;

    execute_phase iDUT_execute (
        .pc_in              (pc_reg),
        .o_rs1_rdata_in     (o_rs1_rdata),
        .o_rs2_rdata_in     (o_rs2_rdata),
        .o_immediate        (o_immediate),
        .jump               (jump),
        .jalr               (jalr),
        .branch             (branch),
        .branch_type        (branch_type),
        .i_opsel            (i_opsel),
        .i_sub              (i_sub),
        .i_unsigned         (i_unsigned),
        .i_arith            (i_arith),
        .auipc              (auipc),
        .i_alu_src          (i_alu_src),
        .pc_out             (pc_next),
        .o_result           (alu_result)
    );

    /////////////////////////////////////
    // Memory Phase
    /////////////////////////////////////
    wire [31:0] load_mux_out;

    memory_phase iDUT_memory (
        .alu_result         (alu_result),
        .load_sel           (load_sel),
        .store_sel          (store_sel),
        .dmem_ren           (dmem_ren),
        .dmem_wen           (dmem_wen),
        .o_rs2_rdata        (o_rs2_rdata),
        .i_dmem_rdata       (i_dmem_rdata),
        .o_dmem_addr        (o_dmem_addr),
        .o_dmem_ren         (o_dmem_ren),
        .o_dmem_wen         (o_dmem_wen),
        .o_dmem_wdata       (o_dmem_wdata),
        .o_dmem_mask        (o_dmem_mask),
        .load_mux_out       (load_mux_out)
    );

    /////////////////////////////////////
    // Writeback Phase
    /////////////////////////////////////
    writeback_phase iDUT_writeback (
        .rd_dest_select     (rd_dest_select),
        .alu_result         (alu_result),
        .pc_plus_4          (pc_plus_4),
        .o_immediate        (o_immediate),
        .load_mux_out       (load_mux_out),
        .writeback_mux_out  (writeback_mux_out)
    );

    /////////////////////////////////////
    // Retire Interface - hart comments
    /////////////////////////////////////
    assign o_retire_valid     = ~i_rst;
    assign o_retire_inst      = instruction;
    assign o_retire_pc        = pc_reg;
    assign o_retire_next_pc   = pc_next;

    assign o_retire_rs1_raddr = instruction[19:15];
    assign o_retire_rs2_raddr = instruction[24:20];
    assign o_retire_rd_waddr  = i_rd_wen ? instruction[11:7] : 5'd0;

    assign o_retire_rs1_rdata = o_rs1_rdata;
    assign o_retire_rs2_rdata = o_rs2_rdata;
    assign o_retire_rd_wdata  = writeback_mux_out;

    // DO NOT FORGOR THIS
    assign o_retire_halt = (instruction == 32'h00100073);

    // Trap on misaligned instruction fetch target or misaligned data access
    wire misaligned_fetch = (jump | jalr | branch) & (pc_next[1:0] != 2'b00);
    wire misaligned_dmem  = (dmem_wen & (store_sel == 3'b010) & (alu_result[1:0] != 2'b00)) |
                            (dmem_wen & (store_sel == 3'b001) & (alu_result[0]   != 1'b0))  |
                            (dmem_ren & (load_sel  == 3'b010) & (alu_result[1:0] != 2'b00)) |
                            (dmem_ren & (load_sel  == 3'b001) & (alu_result[0]   != 1'b0));
    assign o_retire_trap  = misaligned_fetch | misaligned_dmem;

endmodule

`default_nettype wire

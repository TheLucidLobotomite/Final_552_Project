module IDtoEX (
    
);

endmodule
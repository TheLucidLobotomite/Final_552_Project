module moduleName (
    
) (
    ports
);
    
endmodule